module ldr_writeback_unit(
    // pipeline unit ports
    input clk,
    input rst_n,
    input [31:0] instr_in,
    // controller signals
    output w_en_ldr
);

// pipeline unit ports
wire [6:0] opcode_decoded;

// controller ports
reg w_en_ldr_reg;
assign w_en_ldr = w_en_ldr_reg;

// pipeline unit module
writeback_pipeline_unit writeback_pipeline_unit(
    .clk(clk),
    .rst_n(rst_n),
    .instr_in(instr_in),
    .opcode(opcode_decoded)
);

// controller module
always_comb begin
    // default values
    w_en_ldr_reg = 1'b0;

    if (opcode_decoded[6:4] == 3'b110 || opcode_decoded[6:3] == 4'b1000) begin
        //w_en_ldr_reg
        w_en_ldr_reg = 1'b1;
    end
end
endmodule: ldr_writeback_unit