module fetch_wait_unit();
    // does nothing
endmodule: fetch_wait_unit