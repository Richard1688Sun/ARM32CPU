module ldr_writeback_unit();
endmodule: ldr_writeback_unit