module fetch_unit();
// does nothing
endmodule: fetch_unit