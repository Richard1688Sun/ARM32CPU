module memory_wait_unit();
endmodule: memory_wait_unit