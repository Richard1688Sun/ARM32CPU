module memory_unit();
endmodule: memory_unit